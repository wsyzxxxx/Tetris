module vga_controller(iRST_n,
                      iVGA_CLK,
                      oBLANK_n,
                      oHS,
                      oVS,
                      b_data,
                      g_data,
                      r_data,
							 vga_data,
							 vga_addr,
							 vga_wren,
							 write_clk,
							 block_wren,
							 inscore,
							 enscore);
input iRST_n;
input iVGA_CLK;
input block_wren;
input [7:0] vga_data;
input [18:0] vga_addr;
input write_clk;
input vga_wren;
input [31:0] inscore;
input enscore;
output reg oBLANK_n;
output reg oHS;
output reg oVS;
output [7:0] b_data;
output [7:0] g_data;  
output [7:0] r_data;                        
////////////////////
reg [7:0] block_index;
reg [202:0] block_data;                
reg [18:0] ADDR;
reg [23:0] bgr_data;
wire [7:0] index;
wire [23:0] bgr_data_raw;
wire cBLANK_n,cHS,cVS,rst;
wire qout;
wire VGA_CLK_n;
////
assign rst = ~iRST_n;
video_sync_generator LTM_ins (.vga_clk(iVGA_CLK),
                              .reset(rst),
                              .blank_n(cBLANK_n),
                              .HS(cHS),
                              .VS(cVS));
////
////Addresss generator
always@(posedge iVGA_CLK,negedge iRST_n)
begin
  if (!iRST_n)
     ADDR=19'd0;
  else if (cHS==1'b0 && cVS==1'b0)
     ADDR=19'd0;
  else if (cBLANK_n==1'b1) begin
     ADDR=ADDR+19'd1;
  end
end
always@(posedge VGA_CLK_n) begin
  block_data[block_index] = qout;
  if (block_index == 8'd202)
	  block_index = 8'd0;
  else
     block_index = block_index + 8'd1;
end
//////////////////////////
blocks blocks_ram_inst (
	.data (vga_data[0]),
	.rdaddress (block_index),
	.rdclock (VGA_CLK_n),
	.wraddress (vga_addr[7:0]),
	.wrclock (write_clk),
	.wren (block_wren),
	.q (qout)
);
//////INDEX addr.
assign VGA_CLK_n = ~iVGA_CLK;
img_ram img_ram_inst (
	.data (vga_data),
	.rdaddress (ADDR),
	.rdclock (VGA_CLK_n),
	.wraddress (vga_addr),
	.wrclock (write_clk),
	.wren (vga_wren),
	.q (index)
);

scoreLatch scoreLatch_inst(
	.d(inscore), 
	.q(oscore),
	.reset(iRST_n), 
	.wren(enscore), 
	.clk(write_clk)
);
//////Add switch-input logic here
wire [7:0] fakeindex;
parameter reg [7:0] oneblock [0:399] = '{8'h2f,8'h2f,8'h20,8'h2a,8'h2e,8'h33,8'h2a,8'h2a,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h23,8'h2f,8'h34,8'h2f,8'h2f,8'h23,8'h31,8'h26,8'h2d,8'h26,8'h20,8'h2c,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h28,8'h2a,8'h29,8'h2e,8'h20,8'h31,8'h20,8'h22,8'h2a,8'h26,8'h28,8'h23,8'h23,8'h23,8'h23,8'h23,8'h23,8'h23,8'h23,8'h23,8'h28,8'h24,8'h22,8'h2b,8'h28,8'h26,8'h28,8'h30,8'h36,8'h35,8'h36,8'h35,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h30,8'h28,8'h2b,8'h31,8'h2e,8'h2d,8'h2a,8'h36,8'h35,8'h36,8'h32,8'h32,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h25,8'h23,8'h24,8'h26,8'h33,8'h26,8'h26,8'h35,8'h36,8'h25,8'h36,8'h32,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h23,8'h2a,8'h27,8'h2a,8'h20,8'h28,8'h36,8'h32,8'h36,8'h25,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h24,8'h26,8'h29,8'h2a,8'h2c,8'h23,8'h35,8'h32,8'h32,8'h36,8'h25,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h32,8'h28,8'h2e,8'h31,8'h26,8'h23,8'h23,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h23,8'h2a,8'h26,8'h26,8'h23,8'h23,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h23,8'h2a,8'h26,8'h26,8'h23,8'h23,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h23,8'h2a,8'h26,8'h26,8'h23,8'h23,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h23,8'h2a,8'h26,8'h26,8'h23,8'h23,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h23,8'h2a,8'h26,8'h26,8'h23,8'h23,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h23,8'h2a,8'h26,8'h26,8'h23,8'h23,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h23,8'h2a,8'h26,8'h26,8'h23,8'h23,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h35,8'h23,8'h2a,8'h26,8'h23,8'h28,8'h28,8'h30,8'h25,8'h36,8'h35,8'h32,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h36,8'h2f,8'h24,8'h34,8'h2f,8'h2a,8'h24,8'h28,8'h23,8'h23,8'h24,8'h28,8'h23,8'h23,8'h23,8'h23,8'h23,8'h23,8'h23,8'h23,8'h2f,8'h2b,8'h37,8'h26,8'h34,8'h29,8'h22,8'h2b,8'h24,8'h2a,8'h26,8'h2e,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h2a,8'h24,8'h37,8'h26,8'h28,8'h2f,8'h2e,8'h2b,8'h31,8'h26,8'h27,8'h2b,8'h31,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h26,8'h34,8'h26,8'h28,8'h2f};
parameter reg [7:0] zero [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h54, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h54, 8'h55, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] one [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] two [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h55, 8'h54, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] three [0:509] ='{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4d, 8'h54, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h55, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] four [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] five [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] six [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h4f, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h54, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] seven [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] eight [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h55, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h54, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h55, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h54, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] nine [0:509] = '{8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h54, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h55, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4f, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h43, 8'h43, 8'h43, 8'h43, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h54, 8'h4f, 8'h55, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h43, 8'h43, 8'h43, 8'h43, 8'h55, 8'h4f, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d, 8'h4d};
parameter reg [7:0] over [0:19999] = '{8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5e, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5e, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h5b, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h5e, 8'h5e, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5e, 8'h59, 8'h5c, 8'h5e, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5b, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5e, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h5b, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h5b, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h5e, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h59, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5e, 8'h5b, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5e, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h5e, 8'h59, 8'h5e, 8'h5c, 8'h5e, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5b, 8'h5e, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5c, 8'h59, 8'h5c, 8'h5e, 8'h5c, 8'h59, 8'h5e, 8'h5c, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59};
parameter reg [7:0] welcome [0:19999] = '{8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5d, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5d, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5f, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5f, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5f, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5f, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5f, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5b, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h59, 8'h59, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h5d, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5d, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5a, 8'h5f, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5f, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h5b, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h5f, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5b, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h5f, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h5b, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h58, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5b, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5b, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h5b, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5f, 8'h5a, 8'h5f, 8'h5b, 8'h5a, 8'h5f, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h60, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5d, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5b, 8'h59, 8'h59, 8'h5d, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5b, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h59, 8'h5b, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5f, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h5d, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h5d, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h5d, 8'h5d, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5b, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5d, 8'h59, 8'h5f, 8'h59, 8'h59, 8'h58, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h60, 8'h60, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h5a, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5d, 8'h60, 8'h60, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5f, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h5f, 8'h58, 8'h5a, 8'h60, 8'h59, 8'h5f, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5d, 8'h59, 8'h5f, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h58, 8'h5a, 8'h5b, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h58, 8'h59, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5d, 8'h5d, 8'h5b, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5d, 8'h5d, 8'h5a, 8'h5b, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5a, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5b, 8'h5d, 8'h5b, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h59, 8'h5d, 8'h60, 8'h5d, 8'h5d, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h60, 8'h60, 8'h60, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5d, 8'h5a, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5b, 8'h5a, 8'h60, 8'h5d, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h5b, 8'h5d, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h5a, 8'h5f, 8'h60, 8'h5f, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h5a, 8'h5d, 8'h5f, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h5d, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h5d, 8'h5f, 8'h5f, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5d, 8'h5f, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5d, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5d, 8'h58, 8'h5a, 8'h60, 8'h60, 8'h5d, 8'h59, 8'h5a, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h5a, 8'h5a, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5f, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5d, 8'h5b, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5b, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5f, 8'h5f, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5d, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h5f, 8'h5d, 8'h5d, 8'h5b, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5b, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h59, 8'h5d, 8'h5d, 8'h5a, 8'h5b, 8'h59, 8'h5b, 8'h5a, 8'h58, 8'h5a, 8'h5b, 8'h5d, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5b, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5b, 8'h59, 8'h5b, 8'h5b, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5d, 8'h5b, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5b, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h5d, 8'h5b, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h5d, 8'h5d, 8'h5d, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5f, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h58, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5f, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h59, 8'h59, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5f, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5d, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h5f, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5b, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5b, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5f, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h5b, 8'h5b, 8'h5f, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5f, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5f, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h5a, 8'h5f, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5d, 8'h59, 8'h5f, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5f, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h59, 8'h59, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5d, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h58, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h59, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h59, 8'h5b, 8'h59, 8'h5b, 8'h5b, 8'h5b, 8'h59, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h5b, 8'h5d, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5f, 8'h59, 8'h5b, 8'h5b, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5d, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5a, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5f, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h59, 8'h5d, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5d, 8'h59, 8'h5f, 8'h5b, 8'h5b, 8'h5d, 8'h5d, 8'h60, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5d, 8'h5d, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h5d, 8'h5d, 8'h5d, 8'h5d, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5b, 8'h5b, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h59, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5d, 8'h5d, 8'h59, 8'h59, 8'h59, 8'h5b, 8'h5d, 8'h5a, 8'h5a, 8'h60, 8'h59, 8'h5b, 8'h60, 8'h60, 8'h5a, 8'h5d, 8'h5b, 8'h5d, 8'h60, 8'h60, 8'h5a, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5d, 8'h59, 8'h59, 8'h5d, 8'h60, 8'h5a, 8'h60, 8'h59, 8'h59, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5f, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h60, 8'h5a, 8'h5a, 8'h5f, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h58, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5f, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5f, 8'h5f, 8'h5f, 8'h5a, 8'h5a, 8'h5f, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h58, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h60, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5f, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h5a, 8'h60, 8'h60, 8'h5a, 8'h5a, 8'h60, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a, 8'h5a};
parameter reg [7:0] pause [0:19999] = '{8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h63, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h63, 8'h63, 8'h64, 8'h63, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h62, 8'h63, 8'h63, 8'h65, 8'h65, 8'h62, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h64, 8'h65, 8'h65, 8'h62, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h62, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h64, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h62, 8'h63, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h63, 8'h63, 8'h64, 8'h63, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h64, 8'h63, 8'h63, 8'h63, 8'h63, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h62, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h65, 8'h63, 8'h64, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h63, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h62, 8'h65, 8'h62, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h62, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h63, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h62, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h64, 8'h65, 8'h65, 8'h63, 8'h65, 8'h65, 8'h65, 8'h62, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h62, 8'h65, 8'h64, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h63, 8'h63, 8'h64, 8'h63, 8'h63, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h64, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h64, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h65, 8'h65, 8'h63, 8'h64, 8'h63, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h64, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h63, 8'h63, 8'h63, 8'h63, 8'h63, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h61, 8'h64, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h65, 8'h61, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h65, 8'h61, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h64, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h64, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h64, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h62, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h61, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h61, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h61, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h61, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h61, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h65, 8'h62, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h62, 8'h65, 8'h62, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65, 8'h65};
integer x, y;
integer actualX, actualY, relativeX, relativeY, xInside, yInside;
localparam upboader = 40;
localparam downboader = 440;
localparam leftboader = 100;
localparam rightboader = 300;
localparam scoreUp = 90;
localparam scoreDown = 120;
localparam scoreLeft = 460;
localparam scoreRight = 562;
reg [7:0] input_index;
wire [20:0] score;
wire [31:0] oscore;

assign score = oscore[20:0];

always@(negedge VGA_CLK_n) begin
	actualX = ADDR % 19'd640;
	actualY = ADDR / 19'd640;
	if (actualX >= leftboader && actualX < rightboader && actualY >= upboader && actualY < downboader) begin
		xInside = (actualX - leftboader) % 20;
		yInside = (actualY - upboader) % 20;
		relativeX = (actualX - leftboader) / 20 + 2;
		relativeY = (actualY - upboader) / 20;
		input_index = block_data[relativeX + relativeY*10] ? oneblock[xInside + yInside * 20] /*fakebg[ADDR]*/ : index;
	end else if (actualX >= scoreLeft && actualX < scoreRight && actualY >= scoreUp && actualY < scoreDown) begin
		relativeX = (actualX - scoreLeft) / 17;
		xInside = (actualX - scoreLeft) % 17;
		yInside = actualY - scoreUp;
		if (relativeX == 0) begin
			case ((score / 19'd100000) % 10) 
			30'd0: begin
				input_index = zero[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd1: begin
				input_index = one[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd2: begin
				input_index = two[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd3: begin
				input_index = three[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd4: begin
				input_index = four[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd5: begin
				input_index = five[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd6: begin
				input_index = six[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd7: begin
				input_index = seven[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd8: begin
				input_index = eight[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd9: begin
				input_index = nine[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			default: begin
				input_index = index;
			end
			endcase
		end else if (relativeX == 1) begin
			case ((score / 19'd10000) % 10) 
			30'd0: begin
				input_index = zero[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd1: begin
				input_index = one[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd2: begin
				input_index = two[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd3: begin
				input_index = three[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd4: begin
				input_index = four[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd5: begin
				input_index = five[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd6: begin
				input_index = six[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd7: begin
				input_index = seven[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd8: begin
				input_index = eight[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd9: begin
				input_index = nine[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			default: begin
				input_index = index;
			end
			endcase
		end else if (relativeX == 2) begin
			case ((score / 19'd1000) % 10) 
			30'd0: begin
				input_index = zero[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd1: begin
				input_index = one[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd2: begin
				input_index = two[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd3: begin
				input_index = three[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd4: begin
				input_index = four[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd5: begin
				input_index = five[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd6: begin
				input_index = six[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd7: begin
				input_index = seven[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd8: begin
				input_index = eight[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd9: begin
				input_index = nine[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			default: begin
				input_index = index;
			end
			endcase
		end else if (relativeX == 3) begin
			case ((score / 19'd100) % 10) 
			30'd0: begin
				input_index = zero[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd1: begin
				input_index = one[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd2: begin
				input_index = two[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd3: begin
				input_index = three[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd4: begin
				input_index = four[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd5: begin
				input_index = five[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd6: begin
				input_index = six[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd7: begin
				input_index = seven[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd8: begin
				input_index = eight[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd9: begin
				input_index = nine[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			default: begin
				input_index = index;
			end
			endcase
		end else if (relativeX == 4) begin
			case ((score / 19'd10) % 10) 
			30'd0: begin
				input_index = zero[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd1: begin
				input_index = one[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd2: begin
				input_index = two[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd3: begin
				input_index = three[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd4: begin
				input_index = four[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd5: begin
				input_index = five[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd6: begin
				input_index = six[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd7: begin
				input_index = seven[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd8: begin
				input_index = eight[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd9: begin
				input_index = nine[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			default: begin
				input_index = index;
			end
			endcase
		end else if (relativeX == 5) begin
			case (score % 10) 
			30'd0: begin
				input_index = zero[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd1: begin
				input_index = one[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd2: begin
				input_index = two[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd3: begin
				input_index = three[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd4: begin
				input_index = four[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd5: begin
				input_index = five[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd6: begin
				input_index = six[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd7: begin
				input_index = seven[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd8: begin
				input_index = eight[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			30'd9: begin
				input_index = nine[xInside + yInside*17] == 8'h4d ? index : 8'h43;
			end
			default: begin
				input_index = index;
			end
			endcase
		end
	end else begin
		input_index = index;
	end
	if (oscore[30]) begin
		if (actualX >= 220 && actualX < 420 && actualY >= 190 && actualY < 290) begin
			input_index = welcome[actualX - 220 + (actualY - 190) * 200];
		end else begin
			input_index = 8'd96;
		end
	end else if (oscore[29]) begin
		if (actualX >= 220 && actualX < 420 && actualY >= 190 && actualY < 290) begin
			input_index = over[actualX - 220 + (actualY - 190) * 200];
		end
	end else if (oscore[28]) begin
		if (actualX >= 220 && actualX < 420 && actualY >= 190 && actualY < 290) begin
			input_index = pause[actualX - 220 + (actualY - 190) * 200];
		end
	end
end
//////Color table output
img_index	img_index_inst (
	.address ( input_index ),
	.clock ( iVGA_CLK ),
	.q ( bgr_data_raw)
	);	
//////
//////latch valid data at falling edge;
always@(posedge VGA_CLK_n) 
	bgr_data <= bgr_data_raw;
assign b_data = bgr_data[23:16];
assign g_data = bgr_data[15:8];
assign r_data = bgr_data[7:0]; 
///////////////////
//////Delay the iHD, iVD,iDEN for one clock cycle;
always@(negedge iVGA_CLK)
begin
  oHS<=cHS;
  oVS<=cVS;
  oBLANK_n<=cBLANK_n;
end

endmodule
 	















