module Tetris(clock, reset);
    //interface
    input clock;
    input reset;
endmodule
